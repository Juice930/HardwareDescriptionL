LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY REG IS
PORT(RX,BAUD:IN STD_LOGIC;
     RG:OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE REG OF REG IS
BEGIN
	PROCESS(BAUD)
	BEGIN
		IF RISING_EDGE(BAUD) THEN
			RG<=RX;
		END IF;
	END PROCESS;
END REG;