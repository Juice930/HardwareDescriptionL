LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CONTADOR IS 
PORT(BAUD,AVISO_RX:IN STD_LOGIC;
     FIN_CONT8BITS:OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE CONTADOR OF CONTADOR IS
SIGNAL CONTEO:INTEGER RANGE 0 TO 8;
BEGIN
	PROCESS(BAUD)
	BEGIN
		IF AVISO_RX='0' THEN
			FIN_CONT8BITS<='0';
			CONTEO<=0;  
		ELSIF RISING_EDGE(BAUD) THEN
			IF CONTEO=6 THEN
				FIN_CONT8BITS<='1';
			ELSE
				CONTEO<=CONTEO+1;
				FIN_CONT8BITS<='0';
			END IF;
		END IF;
	END PROCESS;
END CONTADOR;