library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity SumRes is

end;

architecture Holi of SumRes is
begin

end Holi;

