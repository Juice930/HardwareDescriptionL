LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY REGRX IS
PORT(BAUD,DESP,RG:IN STD_LOGIC;
     DATOS_RX:BUFFER std_logic_vector(7 downto 0));
END ENTITY;

ARCHITECTURE REGRX OF REGRX IS
BEGIN
	
	PROCESS(BAUD,DESP)
	BEGIN
		IF RISING_EDGE(BAUD) AND DESP='1' THEN
			DATOS_RX(0)<=RG;
			FOR i IN DATOS_RX'length-1 DOWNTO 1 LOOP
				DATOS_RX(i)<=DATOS_RX(i-1);
			END LOOP;
		END IF;
	END PROCESS;
END REGRX;