LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;
ENTITY ADAT IS
PORT (MOTOR,OSC:IN STD_LOGIC;
      INCLINA:IN INTEGER RANGE -3 TO 3;
      SEC:BUFFER INTEGER RANGE 1 TO 8);
END ENTITY;

ARCHITECTURE ADAT OF ADAT IS
SIGNAL CUENTA:INTEGER RANGE 0 TO 24999994;
SIGNAL CLK:STD_LOGIC;
SIGNAL INCLI:INTEGER RANGE -3 TO 3;
BEGIN
  
  PROCESS(OSC)
  BEGIN
  IF MOTOR='1' THEN
  INCLI<=INCLINA;
  END IF;
  IF RISING_EDGE(OSC) THEN
   IF INCLI=-3 OR INCLI=3 THEN
    IF CUENTA=0 THEN
    CUENTA<=1;
    CLK<=NOT CLK;
    ELSE
    CUENTA<=CUENTA-1;
    END IF;
   ELSIF INCLI=-2 OR INCLI=2 THEN
    IF CUENTA=0 THEN
    CUENTA<=2;
    CLK<=NOT CLK;
    ELSE
    CUENTA<=CUENTA-1;
    END IF;
   ELSE
    IF CUENTA=0 THEN
    CUENTA<=4;
    CLK<=NOT CLK;
    ELSE
    CUENTA<=CUENTA-1;
    END IF;
   END IF;
  END IF;
  END PROCESS;  
  
  PROCESS(CLK)
  BEGIN
  IF RISING_EDGE(CLK)THEN
   IF INCLI=3 OR INCLI=2 OR INCLI=1 THEN
   CASE SEC IS
   WHEN 1=>SEC<=2;
   WHEN 2=>SEC<=4;
   WHEN 4=>SEC<=8;
   WHEN 8=>SEC<=1;
   WHEN OTHERS=>SEC<=1;
   END CASE;
   ELSIF INCLI=-1 OR INCLI=-2 OR INCLI=-3 THEN
   CASE SEC IS
   WHEN 8=>SEC<=4;
   WHEN 4=>SEC<=2;
   WHEN 2=>SEC<=1;
   WHEN 1=>SEC<=8;
   WHEN OTHERS=>SEC<=1;
   END CASE;
   ELSE
   SEC<=SEC;
   END IF;
  END IF;
  END PROCESS;

END ADAT;